module testAdd(
 input [63:0] x,
 input [63:0] y,
 input [63:0] z
 );

 assign z = x + y;
 
endmodule
  