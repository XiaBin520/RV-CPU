
import "DPI-C" function void reg_value(input int a, input longint b);

module testBox(
  input  [63:0]  reg_data_0,
  input  [63:0]  reg_data_1,
  input  [63:0]  reg_data_2,
  input  [63:0]  reg_data_3,
  input  [63:0]  reg_data_4,
  input  [63:0]  reg_data_5,
  input  [63:0]  reg_data_6,
  input  [63:0]  reg_data_7,
  input  [63:0]  reg_data_8,
  input  [63:0]  reg_data_9,
  input  [63:0]  reg_data_10,
  input  [63:0]  reg_data_11,
  input  [63:0]  reg_data_12,
  input  [63:0]  reg_data_13,
  input  [63:0]  reg_data_14,
  input  [63:0]  reg_data_15,
  input  [63:0]  reg_data_16,
  input  [63:0]  reg_data_17,
  input  [63:0]  reg_data_18,
  input  [63:0]  reg_data_19,
  input  [63:0]  reg_data_20,
  input  [63:0]  reg_data_21,
  input  [63:0]  reg_data_22,
  input  [63:0]  reg_data_23,
  input  [63:0]  reg_data_24,
  input  [63:0]  reg_data_25,
  input  [63:0]  reg_data_26,
  input  [63:0]  reg_data_27,
  input  [63:0]  reg_data_28,
  input  [63:0]  reg_data_29,
  input  [63:0]  reg_data_30,
  input  [63:0]  reg_data_31
);
 always @(*) begin
   reg_value(0, reg_data_0);
   reg_value(1, reg_data_1);
   reg_value(2, reg_data_2);
   reg_value(3, reg_data_3);
   reg_value(4, reg_data_4);
   reg_value(5, reg_data_5);
   reg_value(6, reg_data_6);
   reg_value(7, reg_data_7);
   reg_value(8, reg_data_8);
   reg_value(9, reg_data_9);
   reg_value(10, reg_data_10);
   reg_value(11, reg_data_11);
   reg_value(12, reg_data_12);
   reg_value(13, reg_data_13);
   reg_value(14, reg_data_14);
   reg_value(15, reg_data_15);
   reg_value(16, reg_data_16);
   reg_value(17, reg_data_17);
   reg_value(18, reg_data_18);
   reg_value(19, reg_data_19);
   reg_value(20, reg_data_20);
   reg_value(21, reg_data_21);
   reg_value(22, reg_data_22);
   reg_value(23, reg_data_23);
   reg_value(24, reg_data_24);
   reg_value(25, reg_data_25);
   reg_value(26, reg_data_26);
   reg_value(27, reg_data_27);
   reg_value(28, reg_data_28);
   reg_value(29, reg_data_29);
   reg_value(30, reg_data_30);
   reg_value(31, reg_data_31);
 end
endmodule
  

    // input  [63:0]  reg_data_0,
    // input  [63:0]  reg_data_1,
    // input  [63:0]  reg_data_2,
    // input  [63:0]  reg_data_3,
    // input  [63:0]  reg_data_4,
    // input  [63:0]  reg_data_5,
    // input  [63:0]  reg_data_6,
    // input  [63:0]  reg_data_7,
    // input  [63:0]  reg_data_8,
    // input  [63:0]  reg_data_9,
    // input  [63:0]  reg_data_10,
    // input  [63:0]  reg_data_11,
    // input  [63:0]  reg_data_12,
    // input  [63:0]  reg_data_13,
    // input  [63:0]  reg_data_14,
    // input  [63:0]  reg_data_15,
    // input  [63:0]  reg_data_16,
    // input  [63:0]  reg_data_17,
    // input  [63:0]  reg_data_18,
    // input  [63:0]  reg_data_19,
    // input  [63:0]  reg_data_20,
    // input  [63:0]  reg_data_21,
    // input  [63:0]  reg_data_22,
    // input  [63:0]  reg_data_23,
    // input  [63:0]  reg_data_24,
    // input  [63:0]  reg_data_25,
    // input  [63:0]  reg_data_26,
    // input  [63:0]  reg_data_27,
    // input  [63:0]  reg_data_28,
    // input  [63:0]  reg_data_29,
    // input  [63:0]  reg_data_30,
    // input  [63:0]  reg_data_31
  